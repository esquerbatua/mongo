module bson

// https://github.com/mongodb/specifications/tree/master/source/bson-corpus/tests
fn test_bson() {

}